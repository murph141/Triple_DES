// $Id: $
// File name:   roundkey.sv
// Created:     3/26/2015
// Author:      Seth Bontrager
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Round Key Generation
