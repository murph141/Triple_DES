// $Id: $
// File name:   io_controller.sv
// Created:     4/1/2015
// Author:      Isaac Sheeley
// Lab Section: 4
// Version:     1.0  Initial Design Entry
// Description: io controller
