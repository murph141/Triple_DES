// $Id: $
// File name:   PBox.sv
// Created:     4/1/2015
// Author:      Anthony Kang
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Permutation Box
module PBox(
  input wire [32:0] data,
  output wire [32:0] p_data
);