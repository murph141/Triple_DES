// $Id: $
// File name:   keyExpansion.sv
// Created:     3/26/2015
// Author:      Isaac Sheeley
// Lab Section: 4
// Version:     1.0  Initial Design Entry
// Description: Key expansion algorithm
